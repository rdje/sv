`include "uvm_macros.svh"
`include "class_macros.svh"

package agent_pkg;
  import uvm_pkg::*;
  
  `include "base_agent.svh"
  `include "agent_helper.svh"
  
endpackage : agent_pkg