package uvm_string_pkg;
import uvm_pkg::*;

typedef string sa_t[$];

`include "uvm_string.svh"
`include "uvm_string_helper.svh"

endpackage : uvm_string_pkg 