package reg_pkg;
import uvm_pkg::*;

`include "base_reg.svh"
`include "base_reg_field.svh"

endpackage : reg_pkg