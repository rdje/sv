class base_reg  extends uvm_reg;
`uvm_object_utils(base_reg)

typedef base_reg this_type;

// Function: new
//
function new();
  
endfunction : new

// Function: write_reg
// Function: read_reg
// Function: update_reg

endclass : base_reg