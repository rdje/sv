
`include "class_macros.svh"

package sb_pkg;
uvm_pkg::*;
event_pkg::*;
  
`include "base_scoreboard.svh"

endpackge : sb_pkg