`include "uvm_macros.svh"
`include "class_macros.svh"

package env_pkg;
  import uvm_pkg::*;
  
  `include "base_env.svh"
  `include "env_helper.svh"
  
endpackage : env_pkg